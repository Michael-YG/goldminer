`ifndef __SHA256_INCL_SVH__
`define __SHA256_INCL_SVH__

`define SHA256_H0 32'h6a09e667 
`define SHA256_H1 32'hbb67ae85
`define SHA256_H2 32'h3c6ef372
`define SHA256_H3 32'ha54ff53a
`define SHA256_H4 32'h510e527f
`define SHA256_H5 32'h9b05688c
`define SHA256_H6 32'h1f83d9ab
`define SHA256_H7 32'h5be0cd19

`endif
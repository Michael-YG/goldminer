`ifndef __SHA256_INCL_SVH__
`define __SHA256_INCL_SVH__

`define SHA256_H0 0x6a09e667 
`define SHA256_H1 0xbb67ae85
`define SHA256_H2 0x3c6ef372
`define SHA256_H3 0xa54ff53a
`define SHA256_H4 0x510e527f
`define SHA256_H5 0x9b05688c
`define SHA256_H6 0x1f83d9ab
`define SHA256_H7 0x5be0cd19

`endif